package apb_pkg;
`include "apb_transaction.sv"
`include "apb_genarator.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_scoreboard.sv"
`include "apb_env.sv"
endpackage